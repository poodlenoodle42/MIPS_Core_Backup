`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/12/2021 04:19:35 PM
// Design Name: 
// Module Name: stall_unit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module stall_unit(
    input rf_stall,
    input mult_div_stall,
    input forwarding,
    output stall_cu,
    output stall_rd,
    output reset_rd,
    output stall_ex,
    output stall_rf
    );
    

endmodule
